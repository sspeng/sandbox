netcdf pism_overrides {
    variables:
    byte pism_overrides;

    pism_overrides:sia_enhancement_factor = 3.0;
    pism_overrides:sia_enhancement_factor_doc = "; Flow enhancement factor for SIA";

    pism_overrides:do_pseudo_plastic_till = "yes";
    pism_overrides:do_pseudo_plastic_till_doc = "Use the pseudo-plastic till model.";

    pism_overrides:pseudo_plastic_q = 0.25;
    pism_overrides:pseudo_plastic_q_doc = "; The exponent of the pseudo-plastic basal resistance model";

    pism_overrides:till_pw_fraction = 0.95;
    pism_overrides:till_pw_fraction_doc = "pure number; pore water pressure is this fraction of overburden";

    pism_overrides:epsilon_ssafd = 1.0e13;
    pism_overrides:epsilon_ssafd_doc = "Pa s m;  Initial amount of regularization in computation of product of effective viscosity nu and thickness H, in SSAFD object.  This quantity is increased if the outer (Picard) iteration is not converging.  This default value for nu * H comes e.g. from a hardness (bar B)=1.9e8 Pa s^(1/3) [\\ref MacAyealetal] and a typical strain rate of 0.001 a-1, giving nu = (bar B) / (2 * 0.001^(2/3)) = 9.49e+14 Pa s ~~ 30 MPa yr, the value in [\\ref Ritzetal2001], and a thickness of H = 10.5 m.";

    pism_overrides:reference_date = "1989-1-1";
    pism_overrides:reference_date_doc = "year-month-day; reference date used in PISM output files";

    pism_overrides:calendar = "360_day";
    pism_overrides:calendar_doc = "The CF calendar keyword in PISM output files.";

    pism_overrides:institution = "University of Alaska Fairbanks";
    pism_overrides:institution_doc = "Institution name. This string is written to output files as the 'institution' global attribute.";

    pism_overrides:backup_interval = 5.0;
    pism_overrides:backup_interval_doc = "hours; wall-clock time between automatic backups";

}
